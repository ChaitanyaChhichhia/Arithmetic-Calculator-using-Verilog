/**********************************

Name:- Chaitanya Chhichhia (19BEC018
		 Digvijaysingh Chudasama (19BEC029)
		 
**********************************/
module adder_4bit(a,b,cin,s,coutf);

input [3:0]a,b; //a,b are the 4 bit no.s to be added
input cin;      //cin is the 1 bit input carry
output [3:0]s;  //s is the 4bit final result of addition
output coutf;   //coutf is the generated output carry
//reg [3:0]s;
wire [2:0]cout; //generated internal carries

adder_1bit add1(a[0],b[0],cin,s[0],cout[0]);     //cin is the input carry to the add1
adder_1bit add2(a[1],b[1],cout[0],s[1],cout[1]); //output carry generated by the add1 acts as input carry to add2
adder_1bit add3(a[2],b[2],cout[1],s[2],cout[2]); //output carry generated by the add2 acts as input carry to add3
adder_1bit add4(a[3],b[3],cout[2],s[3],coutf);   //output carry generated by the add2 is the final output carry

endmodule